module csr_file(
  input clk,
  input resetn,

  input [11:0] waddr,
  input [31:0] wdata,
  input        wvalid,

  input [11:0] raddr,
  input        ravalid,
  output wire [31:0] rdata
);



endmodule